// soc_system_sys_3.v

// Generated using ACDS version 18.1 625
//`default_nettype none
`timescale 1 ps / 1 ps
module disparity_gen_system #(
    parameter blk_w = 16,
    parameter blk_h = 16,
    parameter search_blk_h = 24,
    parameter search_blk_w = 48,
    parameter third_w = 240,
    parameter third_h = 480,
    parameter center_w = 304,
    parameter blk_size = blk_w * blk_h,
    parameter output_confidence = 0
    ) (
		input  wire         clk_clk,                                               //                                           clk.clk
		input  wire         reset_reset_n,                                    //                                         reset.reset_n
        // Control and data from top level system
        input  wire [7:0]   bit_pix_bram_mod_0_center_rd_readdata,           // bit_pix_bram_mod_0:rd_data_centerright -> blk_match:srch_rd_data
        output wire [15:0]  blk_match_srch_master_address,                   // blk_match:srch_rd_addr -> bit_pix_bram_mod_0:rd_address_centerright
        input  wire [15:0]  blk_match_ctrl_fsm_0_control_srch_addr,          // blk_match_ctrl_fsm_0:srch_addr -> blk_match:srch_start_address
        input  wire [15:0]  blk_match_ctrl_fsm_0_control_blk_index,          // blk_match_ctrl_fsm_0:blk_index -> blk_match:blk_index
        input  wire         blk_match_ctrl_fsm_0_control_start,              // blk_match_ctrl_fsm_0:bm_start -> blk_match:start
        output wire         blk_match_ctrl_fsm_0_control_done,               // blk_match_ctrl_fsm_0:bm_start -> blk_match:start
        input  wire [15:0]  blk_match_ctrl_fsm_0_control_blk_addr,           // blk_match_ctrl_fsm_0:blk_addr -> blk_match:blk_start_address
        input  wire [7:0]   bit_pix_bram_mod_0_rd_readdata,                  // bit_pix_bram_mod_0:rd_data -> blk_match:blk_rd_data
        output wire [15:0]  blk_match_blk_master_address,                    // blk_match:blk_rd_addr -> bit_pix_bram_mod_0:rd_address
		// Stream to visualize disparity
		output wire         min_dist_finder_avalon_streaming_source_valid,   // min_dist_finder_avalon_streaming_source.valid
		output wire [15:0]  min_dist_finder_avalon_streaming_source_data,    //                                              .data
        // Stream to the filtering system
		output wire [15:0]  min_dist_finder_out_conduit_blk_index,           //             min_dist_finder_out_conduit.blk_index
		output wire [7:0]   min_dist_finder_out_conduit_sum,                 //                                              .sum
		output wire [7:0]   confidence,                 //                                              .sum
		output wire [15:0]  min_out_coords,                 //                                              .sum
		output wire [blk_size-1:0]  min_xors,                 //                                              .sum
		output wire min_sum_valid                 //                                              .sum
	);

	wire          hamming_dist_out_conduit_valid;               // hamming_dist:sum_valid -> min_dist_finder:sum_valid
	wire   [15:0] hamming_dist_out_conduit_blk_coords;          // hamming_dist:out_coords -> min_dist_finder:out_coords
	wire   [15:0] hamming_dist_out_conduit_blk_index;           // hamming_dist:blk_index_o -> min_dist_finder:blk_index_o
	wire    [7:0] hamming_dist_out_conduit_sum;                 // hamming_dist:sum -> min_dist_finder:sum
	wire          blk_match_result_conduit_blks_valid;          // blk_match:blks_valid -> hamming_dist:blks_valid
	wire  [blk_size-1:0] blk_match_result_conduit_srch_block;          // blk_match:srch_block -> hamming_dist:left
	wire   [15:0] blk_match_result_conduit_blk_index;           // blk_match:blk_index_o -> hamming_dist:blk_index_i
	wire   [15:0] blk_match_result_conduit_coords_out;          // blk_match:coords_out -> hamming_dist:in_coords
	wire  [blk_size-1:0] blk_match_result_conduit_blk_block;           // blk_match:blk_block -> hamming_dist:right


	block_match_new #(
		.rd_port_w    (8),
		.block_width  (blk_w),
		.block_height (blk_h),
		.search_blk_w (search_blk_w),
		.search_blk_h (search_blk_h),
		.center_w     (center_w),
		.third_w      (third_w)
    ) blk_match (
		.clk                (clk_clk),                                      //          clock.clk
		.reset              (~reset_reset_n),           //          reset.reset
		.blk_index          (blk_match_ctrl_fsm_0_control_blk_index), //   ctrl_conduit.blk_index
		.start              (blk_match_ctrl_fsm_0_control_start),     //               .start
		.done               (blk_match_ctrl_fsm_0_control_done),                                             //               .done
		.blk_start_address  (blk_match_ctrl_fsm_0_control_blk_addr),  //               .blk_addr
		.srch_start_address (blk_match_ctrl_fsm_0_control_srch_addr), //               .srch_addr
		.blk_block          (blk_match_result_conduit_blk_block),     // result_conduit.blk_block
		.blk_index_o        (blk_match_result_conduit_blk_index),     //               .blk_index
		.srch_block         (blk_match_result_conduit_srch_block),    //               .srch_block
		.coords_out         (blk_match_result_conduit_coords_out),    //               .coords_out
		.blks_valid         (blk_match_result_conduit_blks_valid),    //               .blks_valid
		.srch_rd_addr       (blk_match_srch_master_address),          //    srch_master.address
		.srch_rd_data       (bit_pix_bram_mod_0_center_rd_readdata),   //               .readdata
		.blk_rd_addr        (blk_match_blk_master_address),           //     blk_master.address
		.blk_rd_data        (bit_pix_bram_mod_0_rd_readdata)          //               .readdata
	);

    logic [blk_size - 1:0]  hd_xors;

	hamming_dist_new #(
		.blk_size    (blk_size),
		.lut_bits_in (4)
	) hamming_dist (
		.clk         (clk_clk),                                   //       clock.clk
		.reset       (~reset_reset_n),        //       reset.reset
		.blk_index_o (hamming_dist_out_conduit_blk_index),  // out_conduit.blk_index
		.sum_valid   (hamming_dist_out_conduit_valid),      //            .valid
		.sum         (hamming_dist_out_conduit_sum),        //            .sum
		.xors        (hd_xors),                                          //            .xors
		.out_coords  (hamming_dist_out_conduit_blk_coords), //            .blk_coords
		.right       (blk_match_result_conduit_blk_block),  //  in_conduit.blk_block
		.left        (blk_match_result_conduit_srch_block), //            .srch_block
		.blk_index_i (blk_match_result_conduit_blk_index),  //            .blk_index
		.blks_valid  (blk_match_result_conduit_blks_valid), //            .blks_valid
		.in_coords   (blk_match_result_conduit_coords_out)  //            .coords_out
	);
    
	min_dist_finder #(
		.blk_h        (blk_h),
		.blk_w        (blk_w),
        .third_h      (third_h),
		.search_blk_w (search_blk_w),
		.search_blk_h (search_blk_h),
        .output_confidence  (output_confidence)
	) min_dist_finder (
		.clk             (clk_clk),                                             //                   clock.clk
		.reset           (~reset_reset_n),                      //                   reset.reset
        
        .xors            (hd_xors),
		.sum             (hamming_dist_out_conduit_sum),                  //              in_conduit.sum
		.out_coords      (hamming_dist_out_conduit_blk_coords),           //                        .blk_coords
		.sum_valid       (hamming_dist_out_conduit_valid),                //                        .valid
		.blk_index_o     (hamming_dist_out_conduit_blk_index),            //                        .blk_index
        
		.stream_out_valid(min_dist_finder_avalon_streaming_source_valid), // avalon_streaming_source.valid
		.stream_out      (min_dist_finder_avalon_streaming_source_data),   //                        .data
        
		.min_out_coords  (min_out_coords),   //                        .data
		.min_blk_index_o (min_dist_finder_out_conduit_blk_index),         //             out_conduit.blk_index
        .min_xors        (min_xors),
		.min_sum         (min_dist_finder_out_conduit_sum),               //                        .sum
		.min_sumh        (),              //                        .data
		.confidence      (confidence),   //                        .data
        .min_sum_valid   (min_sum_valid)
	);
endmodule
