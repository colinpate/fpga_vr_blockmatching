// soc_system_sys_2.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module bit_pixel_conversion_system #(
    parameter third_cols = 240,
    parameter third_rows = 480,
    parameter center_cols = 304
    ) (
		output wire [15:0]  bram_writer_0_avalon_master_writedata,                 //             bram_writer_0_avalon_master.writedata
		output wire         bram_writer_0_avalon_master_write,                     //                                        .write
		output wire [15:0]  bram_writer_0_avalon_master_address,                   //                                        .address
		output wire [1:0]   bram_writer_0_avalon_master_third,                   //                                        .address
		output wire [15:0]  bram_writer_0_avalon_master_1_writedata,               //           bram_writer_0_avalon_master_1.writedata
		output wire         bram_writer_0_avalon_master_1_write,                   //                                        .write
		output wire [15:0]  bram_writer_0_avalon_master_1_address,                 //                                        .address
		output wire [1:0]   bram_writer_0_avalon_master_1_third,                 //                                        .address
		input  wire         bram_writer_0_bm_status_conduit_bm_idle,               //         bram_writer_0_bm_status_conduit.bm_idle
		input  wire         bram_writer_0_bm_status_conduit_bm_working_buf,        //                                        .bm_working_buf
		output wire [3:0]   bram_writer_0_bm_status_conduit_image_number,          //                                        .image_number
		output wire [3:0]   bram_writer_0_bm_status_conduit_b_image_number,        //       bram_writer_0_bm_status_conduit_b.image_number
		input  wire [1:0]   ddr3_reader_fsm_0_cam_0_ptr_sink_data,                 //        ddr3_reader_fsm_0_cam_0_ptr_sink.data
		output wire         ddr3_reader_fsm_0_cam_0_ptr_sink_ready,                //                                        .ready
		input  wire         ddr3_reader_fsm_0_cam_0_ptr_sink_valid,                //                                        .valid
		input  wire [31:0]  ddr3_reader_fsm_0_cam_0_start_start_addr,              //           ddr3_reader_fsm_0_cam_0_start.start_addr
		input  wire [1:0]   ddr3_reader_fsm_0_cam_1_ptr_sink_data,                 //        ddr3_reader_fsm_0_cam_1_ptr_sink.data
		output wire         ddr3_reader_fsm_0_cam_1_ptr_sink_ready,                //                                        .ready
		input  wire         ddr3_reader_fsm_0_cam_1_ptr_sink_valid,                //                                        .valid
		input  wire [31:0]  ddr3_reader_fsm_0_cam_1_start_start_addr,              //           ddr3_reader_fsm_0_cam_1_start.start_addr
		output wire [26:0]  ddr3_reader_vertical_0_ddr3_read_master_address,       // ddr3_reader_vertical_0_ddr3_read_master.address
		input  wire [255:0] ddr3_reader_vertical_0_ddr3_read_master_readdata,      //                                        .readdata
		output wire         ddr3_reader_vertical_0_ddr3_read_master_read,          //                                        .read
		input  wire         ddr3_reader_vertical_0_ddr3_read_master_waitrequest,   //                                        .waitrequest
		input  wire         ddr3_reader_vertical_0_ddr3_read_master_readdatavalid, //                                        .readdatavalid
		output wire [3:0]   ddr3_reader_vertical_0_ddr3_read_master_burstcount,    //                                        .burstcount
		input  wire         ddr3clk_clk,                                           //                                 ddr3clk.clk
		input  wire         ddr3clk_reset_reset_n,                                 //                           ddr3clk_reset.reset_n
		input  wire         pclk_clk,                                              //                                    pclk.clk
		input  wire         pclk_reset_reset_n                                     //                              pclk_reset.reset_n
	);

	wire          gray_vertical_filter_bank_0_avalon_streaming_source_valid; // gray_vertical_filter_bank_0:bit_pixels_valid -> bram_writer_0:bit_pix_valid
	wire   [23:0] gray_vertical_filter_bank_0_avalon_streaming_source_data;  // gray_vertical_filter_bank_0:bit_pixels -> bram_writer_0:bit_pix
	wire          bram_writer_0_fifo_almost_full_source_data;                // bram_writer_0:fifo_almost_full -> ddr3_reader_vertical_0:pix_fifo_almost_full
	wire          ddr3_reader_vertical_0_pixel_source_valid;                 // ddr3_reader_vertical_0:pixel_valid -> gray_vertical_filter_bank_0:pixel_in_valid
	wire  [263:0] ddr3_reader_vertical_0_pixel_source_data;                  // ddr3_reader_vertical_0:pixel_data -> gray_vertical_filter_bank_0:pixel_in
	wire          ddr3_reader_fsm_0_read_addr_src_valid;                     // ddr3_reader_fsm_0:read_addr_valid -> ddr3_reader_vertical_0:start_valid
	wire   [28:0] ddr3_reader_fsm_0_read_addr_src_data;                      // ddr3_reader_fsm_0:read_addr_data -> ddr3_reader_vertical_0:start_data
	wire          ddr3_reader_fsm_0_read_addr_src_ready;                     // ddr3_reader_vertical_0:start_ready -> ddr3_reader_fsm_0:read_addr_ready
	wire          rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [bram_writer_0:reset, ddr3_reader_vertical_0:pclk_reset, gray_vertical_filter_bank_0:reset]
	wire          rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> ddr3_reader_vertical_0:ddr3clk_reset

	bit_pixel_rotator_bram #(
		.third_cols     (third_cols),
        .center_cols    (center_cols),
		.third_rows     (third_rows),
		.test_mode      (0)
	) bram_writer_0 (
		.clk              (pclk_clk),                                                  //                   clock.clk
		.reset            (~pclk_reset_reset_n),                            //                   reset.reset
		.pix_out          (bram_writer_0_avalon_master_writedata),                     //           avalon_master.writedata
		.pix_out_wren     (bram_writer_0_avalon_master_write),                         //                        .write
		.pix_out_addr     (bram_writer_0_avalon_master_address),                       //                        .address
		.pix_out_third    (bram_writer_0_avalon_master_third),                       //                        .address
		.bit_pix          (gray_vertical_filter_bank_0_avalon_streaming_source_data),  //            bit_pix_sink.data
		.bit_pix_valid    (gray_vertical_filter_bank_0_avalon_streaming_source_valid), //                        .valid
		.fifo_almost_full (bram_writer_0_fifo_almost_full_source_data),                // fifo_almost_full_source.data
		.bm_idle          (bram_writer_0_bm_status_conduit_bm_idle),                   //       bm_status_conduit.bm_idle
		.bm_working_buf   (bram_writer_0_bm_status_conduit_bm_working_buf),            //                        .bm_working_buf
		.image_number     (bram_writer_0_bm_status_conduit_image_number),              //                        .image_number
		.pix_out_b        (bram_writer_0_avalon_master_1_writedata),                   //         avalon_master_1.writedata
		.pix_out_wren_b   (bram_writer_0_avalon_master_1_write),                       //                        .write
		.pix_out_addr_b   (bram_writer_0_avalon_master_1_address),                     //                        .address
		.pix_out_third_b   (bram_writer_0_avalon_master_1_third),                     //                        .address
		.image_number_b   (bram_writer_0_bm_status_conduit_b_image_number)             //     bm_status_conduit_b.image_number
	);

	ddr3_reader_fsm #(
		.test_mode (1),
        .center_w   (center_cols),
        .third_w    (third_cols)
	) ddr3_reader_fsm_0 (
		.clk             (ddr3clk_clk),                              //          clock.clk
		.reset           (~ddr3clk_reset_reset_n),                   //          reset.reset
		.cam_0_ptr_data  (ddr3_reader_fsm_0_cam_0_ptr_sink_data),    // cam_0_ptr_sink.data
		.cam_0_ptr_ready (ddr3_reader_fsm_0_cam_0_ptr_sink_ready),   //               .ready
		.cam_0_ptr_valid (ddr3_reader_fsm_0_cam_0_ptr_sink_valid),   //               .valid
		.cam_1_ptr_data  (ddr3_reader_fsm_0_cam_1_ptr_sink_data),    // cam_1_ptr_sink.data
		.cam_1_ptr_ready (ddr3_reader_fsm_0_cam_1_ptr_sink_ready),   //               .ready
		.cam_1_ptr_valid (ddr3_reader_fsm_0_cam_1_ptr_sink_valid),   //               .valid
		.cam_0_start     (ddr3_reader_fsm_0_cam_0_start_start_addr), //    cam_0_start.start_addr
		.cam_1_start     (ddr3_reader_fsm_0_cam_1_start_start_addr), //    cam_1_start.start_addr
		.read_addr_ready (ddr3_reader_fsm_0_read_addr_src_ready),    //  read_addr_src.ready
		.read_addr_data  (ddr3_reader_fsm_0_read_addr_src_data),     //               .data
		.read_addr_valid (ddr3_reader_fsm_0_read_addr_src_valid)     //               .valid
	);

	ddr3_reader_grayfilter_short #(
		.frame_third_width (third_cols),
		.center_width      (center_cols),
		.frame_lines       (third_rows),
		.frame_full_width  (768)
	) ddr3_reader_vertical_0 (
		.ddr3clk_reset        (~ddr3clk_reset_reset_n),                    //         ddr3clk_reset.reset
		.pclk_reset           (~pclk_reset_reset_n),                        //            pclk_reset.reset
		.pixel_data           (ddr3_reader_vertical_0_pixel_source_data),              //          pixel_source.data
		.pixel_valid          (ddr3_reader_vertical_0_pixel_source_valid),             //                      .valid
		.pix_fifo_almost_full (bram_writer_0_fifo_almost_full_source_data),            // fifo_almost_full_sink.data
		.start_ready          (ddr3_reader_fsm_0_read_addr_src_ready),                 //       start_addr_sink.ready
		.start_valid          (ddr3_reader_fsm_0_read_addr_src_valid),                 //                      .valid
		.start_data           (ddr3_reader_fsm_0_read_addr_src_data),                  //                      .data
		.ddr3_address         (ddr3_reader_vertical_0_ddr3_read_master_address),       //      ddr3_read_master.address
		.ddr3_readdata        (ddr3_reader_vertical_0_ddr3_read_master_readdata),      //                      .readdata
		.ddr3_read            (ddr3_reader_vertical_0_ddr3_read_master_read),          //                      .read
		.ddr3_waitrequest     (ddr3_reader_vertical_0_ddr3_read_master_waitrequest),   //                      .waitrequest
		.ddr3_readdatavalid   (ddr3_reader_vertical_0_ddr3_read_master_readdatavalid), //                      .readdatavalid
		.ddr3_burstcount      (ddr3_reader_vertical_0_ddr3_read_master_burstcount),    //                      .burstcount
		.pclk                 (pclk_clk),                                              //             pclk_sink.clk
		.ddr3clk              (ddr3clk_clk)                                            //          ddr3clk_sink.clk
	);

	gray_vertical_filter_bank #(
		.n_filters   (16),
		.radius      (8),
		.frame_lines (third_rows)
	) gray_vertical_filter_bank_0 (
		.clk              (pclk_clk),                                                  //                   clock.clk
		.reset            (~pclk_reset_reset_n),                            //                   reset.reset
		.bit_pixels       (gray_vertical_filter_bank_0_avalon_streaming_source_data),  // avalon_streaming_source.data
		.bit_pixels_valid (gray_vertical_filter_bank_0_avalon_streaming_source_valid), //                        .valid
		.pixel_in         (ddr3_reader_vertical_0_pixel_source_data),                  //   avalon_streaming_sink.data
		.pixel_in_valid   (ddr3_reader_vertical_0_pixel_source_valid)                  //                        .valid
	);

endmodule
